interface InterFace ();
    logic [7:0] AIF;
    logic [7:0] BIF;
    logic ENIF;
    logic [3:0] ALU_FUNIF;
    logic CLKIF;
    logic RSTIF;
    logic [15:0] ALU_OUTIF;
endinterface
